`timescale 1ns/1ns
`include "define.sv"

module sm_warp_assign (
	input  clk,                                               // input clock for the system
	input  rst_n, 
	
	
);






endmodule