`timescale 1ns/1ns
`include "define.sv"


module GPGPU_top (


);





endmodule
